`timescale 1ns / 1ps
module system
(
	input clk,
	input rst_n,
);

endmodule