/**
 * File name:	control_unit_if.vh
 * Created:	12/22/2021
 * Author:	Weili An
 * Email:	an107@purdue.edu
 * Version:	1.0 Initial Design Entry
 * Description:	Control/decoder unit interface
 */

`ifndef __CONTROL_UNIT_IF_VH__
`define __CONTROL_UNIT_IF_VH__

`include "rv32ima_pkg.svh"

interface control_unit_if;
    import rv32ima_pkg::*;
    
endinterface // control_unit_if

`endif // __CONTROL_UNIT_IF_VH__