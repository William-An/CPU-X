`timescale 1ns/1ns
module tb_system;
	
endmodule